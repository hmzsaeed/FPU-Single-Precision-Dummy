##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Sun May 29 13:40:23 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO user_proj_example
  CLASS BLOCK ;
  SIZE 933.800000 BY 926.160000 ;
  FOREIGN user_proj_example 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.852 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 0.9534 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 4.606 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 120.593 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 643.632 LAYER met3  ;
    ANTENNAGATEAREA 0.852 LAYER met3  ;
    ANTENNAMAXAREACAR 143.514 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 764.261 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.107277 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1.840000 0.000000 1.980000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4082 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 31.815 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.99 LAYER met2  ;
    ANTENNAMAXAREACAR 14.0833 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 68.4318 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.0519192 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 5.200000 0.490000 5.340000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.465000 0.000000 198.605000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.745000 0.000000 66.885000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.375000 0.000000 200.515000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.555000 0.000000 196.695000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.650000 0.000000 194.790000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.740000 0.000000 192.880000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.830000 0.000000 190.970000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.835000 0.000000 127.975000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.925000 0.000000 126.065000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.015000 0.000000 124.155000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.105000 0.000000 122.245000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.195000 0.000000 120.335000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.290000 0.000000 118.430000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.380000 0.000000 116.520000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.470000 0.000000 114.610000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.560000 0.000000 112.700000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.650000 0.000000 110.790000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.745000 0.000000 108.885000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.835000 0.000000 106.975000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.925000 0.000000 105.065000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.015000 0.000000 103.155000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.105000 0.000000 101.245000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.200000 0.000000 99.340000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.290000 0.000000 97.430000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.380000 0.000000 95.520000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470000 0.000000 93.610000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.560000 0.000000 91.700000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.655000 0.000000 89.795000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.745000 0.000000 87.885000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.835000 0.000000 85.975000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.925000 0.000000 84.065000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.015000 0.000000 82.155000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.110000 0.000000 80.250000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.200000 0.000000 78.340000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.290000 0.000000 76.430000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.380000 0.000000 74.520000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.470000 0.000000 72.610000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.565000 0.000000 70.705000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.655000 0.000000 68.795000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.835000 0.000000 64.975000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.925000 0.000000 63.065000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.020000 0.000000 61.160000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.110000 0.000000 59.250000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.200000 0.000000 57.340000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290000 0.000000 55.430000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.380000 0.000000 53.520000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.475000 0.000000 51.615000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.565000 0.000000 49.705000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.655000 0.000000 47.795000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.745000 0.000000 45.885000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.835000 0.000000 43.975000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.930000 0.000000 42.070000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.020000 0.000000 40.160000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.110000 0.000000 38.250000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.200000 0.000000 36.340000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.290000 0.000000 34.430000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.385000 0.000000 32.525000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.475000 0.000000 30.615000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.565000 0.000000 28.705000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.655000 0.000000 26.795000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.745000 0.000000 24.885000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.840000 0.000000 22.980000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.930000 0.000000 21.070000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.020000 0.000000 19.160000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110000 0.000000 17.250000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.200000 0.000000 15.340000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.295000 0.000000 13.435000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.385000 0.000000 11.525000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.475000 0.000000 9.615000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.565000 0.000000 7.705000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.655000 0.000000 5.795000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8005 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.1745 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 3.750000 0.000000 3.890000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8103 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3215 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 188.920000 0.000000 189.060000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 187.010000 0.000000 187.150000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 185.105000 0.000000 185.245000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 183.195000 0.000000 183.335000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 181.285000 0.000000 181.425000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 179.375000 0.000000 179.515000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 177.465000 0.000000 177.605000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 175.560000 0.000000 175.700000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 173.650000 0.000000 173.790000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 171.740000 0.000000 171.880000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 169.830000 0.000000 169.970000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 167.920000 0.000000 168.060000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 166.015000 0.000000 166.155000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 164.105000 0.000000 164.245000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 162.195000 0.000000 162.335000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 160.285000 0.000000 160.425000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 158.375000 0.000000 158.515000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 156.470000 0.000000 156.610000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 154.560000 0.000000 154.700000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 152.650000 0.000000 152.790000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 150.740000 0.000000 150.880000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 148.830000 0.000000 148.970000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 146.925000 0.000000 147.065000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 145.015000 0.000000 145.155000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 143.105000 0.000000 143.245000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 141.195000 0.000000 141.335000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 139.285000 0.000000 139.425000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 137.380000 0.000000 137.520000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 135.470000 0.000000 135.610000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.3705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 133.560000 0.000000 133.700000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 131.650000 0.000000 131.790000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.8201 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 73.423 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.2 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 3.1621 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 129.740000 0.000000 129.880000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.725000 0.000000 444.865000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.820000 0.000000 442.960000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.910000 0.000000 441.050000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.000000 0.000000 439.140000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090000 0.000000 437.230000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.180000 0.000000 435.320000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.275000 0.000000 433.415000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.365000 0.000000 431.505000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.455000 0.000000 429.595000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.545000 0.000000 427.685000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.635000 0.000000 425.775000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.730000 0.000000 423.870000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.820000 0.000000 421.960000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.910000 0.000000 420.050000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.000000 0.000000 418.140000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.090000 0.000000 416.230000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.185000 0.000000 414.325000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.275000 0.000000 412.415000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.365000 0.000000 410.505000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.455000 0.000000 408.595000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.545000 0.000000 406.685000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.640000 0.000000 404.780000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.730000 0.000000 402.870000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.820000 0.000000 400.960000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910000 0.000000 399.050000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.000000 0.000000 397.140000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.095000 0.000000 395.235000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.185000 0.000000 393.325000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.275000 0.000000 391.415000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.365000 0.000000 389.505000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.455000 0.000000 387.595000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.550000 0.000000 385.690000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.640000 0.000000 383.780000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.730000 0.000000 381.870000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.820000 0.000000 379.960000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.910000 0.000000 378.050000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.005000 0.000000 376.145000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.095000 0.000000 374.235000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.185000 0.000000 372.325000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.275000 0.000000 370.415000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.365000 0.000000 368.505000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.460000 0.000000 366.600000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.550000 0.000000 364.690000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.640000 0.000000 362.780000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730000 0.000000 360.870000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.820000 0.000000 358.960000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.915000 0.000000 357.055000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.005000 0.000000 355.145000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.095000 0.000000 353.235000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.185000 0.000000 351.325000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.275000 0.000000 349.415000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.370000 0.000000 347.510000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.460000 0.000000 345.600000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.550000 0.000000 343.690000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.640000 0.000000 341.780000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.730000 0.000000 339.870000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.825000 0.000000 337.965000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.915000 0.000000 336.055000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.005000 0.000000 334.145000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.095000 0.000000 332.235000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.185000 0.000000 330.325000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.280000 0.000000 328.420000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3087 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1.3825 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 18.532 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 99.304 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 125.187 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 670.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 7.1775 LAYER met4  ;
    ANTENNAMAXAREACAR 27.4067 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 141.632 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.230765 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 326.370000 0.000000 326.510000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.5969 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 177.18 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.968 LAYER met2  ;
    ANTENNAMAXAREACAR 20.4837 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 96.4738 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.190854 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 30.7027 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 164.68 LAYER met3  ;
    ANTENNAGATEAREA 2.952 LAYER met3  ;
    ANTENNAMAXAREACAR 30.8843 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 152.26 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.204404 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 345.547 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1849.48 LAYER met4  ;
    ANTENNAGATEAREA 12.462 LAYER met4  ;
    ANTENNAMAXAREACAR 110.031 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 579.801 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 324.460000 0.000000 324.600000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550000 0.000000 322.690000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.640000 0.000000 320.780000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.735000 0.000000 318.875000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.825000 0.000000 316.965000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.915000 0.000000 315.055000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.005000 0.000000 313.145000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.095000 0.000000 311.235000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.190000 0.000000 309.330000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.280000 0.000000 307.420000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.370000 0.000000 305.510000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.460000 0.000000 303.600000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.550000 0.000000 301.690000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.645000 0.000000 299.785000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.735000 0.000000 297.875000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.825000 0.000000 295.965000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.915000 0.000000 294.055000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.005000 0.000000 292.145000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.100000 0.000000 290.240000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.190000 0.000000 288.330000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.280000 0.000000 286.420000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370000 0.000000 284.510000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.460000 0.000000 282.600000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.555000 0.000000 280.695000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.645000 0.000000 278.785000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.735000 0.000000 276.875000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.825000 0.000000 274.965000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.915000 0.000000 273.055000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.010000 0.000000 271.150000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.100000 0.000000 269.240000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.190000 0.000000 267.330000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.280000 0.000000 265.420000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.370000 0.000000 263.510000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.465000 0.000000 261.605000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.555000 0.000000 259.695000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.645000 0.000000 257.785000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.735000 0.000000 255.875000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.825000 0.000000 253.965000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.920000 0.000000 252.060000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.010000 0.000000 250.150000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.100000 0.000000 248.240000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190000 0.000000 246.330000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.280000 0.000000 244.420000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.375000 0.000000 242.515000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.465000 0.000000 240.605000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.555000 0.000000 238.695000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.645000 0.000000 236.785000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.735000 0.000000 234.875000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.830000 0.000000 232.970000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.920000 0.000000 231.060000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.010000 0.000000 229.150000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.100000 0.000000 227.240000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.190000 0.000000 225.330000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.285000 0.000000 223.425000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.375000 0.000000 221.515000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.465000 0.000000 219.605000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.555000 0.000000 217.695000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.645000 0.000000 215.785000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.740000 0.000000 213.880000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.830000 0.000000 211.970000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.920000 0.000000 210.060000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010000 0.000000 208.150000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.100000 0.000000 206.240000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2259 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7855 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met2  ;
    ANTENNAMAXAREACAR 15.2915 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 58.1572 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.32327 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 204.195000 0.000000 204.335000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.285000 0.000000 202.425000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6038 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.891 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 689.080000 0.000000 689.220000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 687.170000 0.000000 687.310000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 685.260000 0.000000 685.400000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 683.350000 0.000000 683.490000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 681.445000 0.000000 681.585000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 679.535000 0.000000 679.675000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 677.625000 0.000000 677.765000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 675.715000 0.000000 675.855000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 673.805000 0.000000 673.945000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 671.900000 0.000000 672.040000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 669.990000 0.000000 670.130000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 668.080000 0.000000 668.220000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 666.170000 0.000000 666.310000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 664.260000 0.000000 664.400000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 662.355000 0.000000 662.495000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 660.445000 0.000000 660.585000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 658.535000 0.000000 658.675000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 656.625000 0.000000 656.765000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 654.715000 0.000000 654.855000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 652.810000 0.000000 652.950000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 650.900000 0.000000 651.040000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 648.990000 0.000000 649.130000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 647.080000 0.000000 647.220000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 645.170000 0.000000 645.310000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 643.265000 0.000000 643.405000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 641.355000 0.000000 641.495000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 639.445000 0.000000 639.585000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 637.535000 0.000000 637.675000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 635.625000 0.000000 635.765000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 633.720000 0.000000 633.860000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 631.810000 0.000000 631.950000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 629.900000 0.000000 630.040000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 627.990000 0.000000 628.130000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 626.080000 0.000000 626.220000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 624.175000 0.000000 624.315000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 622.265000 0.000000 622.405000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 620.355000 0.000000 620.495000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 618.445000 0.000000 618.585000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 616.535000 0.000000 616.675000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 614.630000 0.000000 614.770000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 612.720000 0.000000 612.860000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 610.810000 0.000000 610.950000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 608.900000 0.000000 609.040000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 606.990000 0.000000 607.130000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 605.085000 0.000000 605.225000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 603.175000 0.000000 603.315000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 601.265000 0.000000 601.405000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 599.355000 0.000000 599.495000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 597.445000 0.000000 597.585000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 595.540000 0.000000 595.680000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 593.630000 0.000000 593.770000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 591.720000 0.000000 591.860000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 589.810000 0.000000 589.950000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 587.900000 0.000000 588.040000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 585.995000 0.000000 586.135000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 584.085000 0.000000 584.225000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 582.175000 0.000000 582.315000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 580.265000 0.000000 580.405000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 578.355000 0.000000 578.495000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 576.450000 0.000000 576.590000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 574.540000 0.000000 574.680000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.94 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 572.630000 0.000000 572.770000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6136 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 107.993 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 570.720000 0.000000 570.860000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.6283 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 108.014 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 568.810000 0.000000 568.950000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5525 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6545 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 566.905000 0.000000 567.045000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.5497 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.6405 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 564.995000 0.000000 565.135000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.6729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2565 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 563.085000 0.000000 563.225000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.158 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 561.175000 0.000000 561.315000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3295 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.5395 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 559.265000 0.000000 559.405000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.158 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 557.360000 0.000000 557.500000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.4235 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 555.450000 0.000000 555.590000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.966 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 553.540000 0.000000 553.680000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.9788 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.786 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 551.630000 0.000000 551.770000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4786 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.285 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 549.720000 0.000000 549.860000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1723 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.7535 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 547.815000 0.000000 547.955000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.87 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 545.905000 0.000000 546.045000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.7764 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.774 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 543.995000 0.000000 544.135000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.9098 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.441 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 542.085000 0.000000 542.225000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.35 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 540.175000 0.000000 540.315000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.3568 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.676 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 538.270000 0.000000 538.410000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.254 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 536.360000 0.000000 536.500000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 4.1628 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 20.706 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 534.450000 0.000000 534.590000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.1534 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 15.659 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 532.540000 0.000000 532.680000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.966 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 530.630000 0.000000 530.770000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.634 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.062 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 528.725000 0.000000 528.865000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.158 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 526.815000 0.000000 526.955000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.35 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 524.905000 0.000000 525.045000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.254 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 522.995000 0.000000 523.135000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.3956 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 16.87 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 521.085000 0.000000 521.225000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.0148 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 14.966 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 519.180000 0.000000 519.320000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.4978 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 17.381 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 517.270000 0.000000 517.410000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.2532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.158 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 515.360000 0.000000 515.500000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.35 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 513.450000 0.000000 513.590000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.8724 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.254 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 511.540000 0.000000 511.680000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 3.8051 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 18.9175 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 509.635000 0.000000 509.775000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.2809 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 1.4916 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.35 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 507.725000 0.000000 507.865000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.983 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4163 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 340.88 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 505.815000 0.000000 505.955000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 503.905000 0.000000 504.045000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 501.995000 0.000000 502.135000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 500.090000 0.000000 500.230000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 498.180000 0.000000 498.320000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 496.270000 0.000000 496.410000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 494.360000 0.000000 494.500000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 492.450000 0.000000 492.590000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 490.545000 0.000000 490.685000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 488.635000 0.000000 488.775000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 486.725000 0.000000 486.865000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 484.815000 0.000000 484.955000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 482.905000 0.000000 483.045000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 481.000000 0.000000 481.140000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 479.090000 0.000000 479.230000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 477.180000 0.000000 477.320000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 475.270000 0.000000 475.410000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 473.360000 0.000000 473.500000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 471.455000 0.000000 471.595000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 469.545000 0.000000 469.685000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 467.635000 0.000000 467.775000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 465.725000 0.000000 465.865000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 463.815000 0.000000 463.955000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 461.910000 0.000000 462.050000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 460.000000 0.000000 460.140000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 458.090000 0.000000 458.230000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 456.180000 0.000000 456.320000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 454.270000 0.000000 454.410000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.397 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 452.365000 0.000000 452.505000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.0845 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 70.944 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 350.997 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.261578 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 450.455000 0.000000 450.595000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4536 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 67.032 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4662 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 341.13 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 448.545000 0.000000 448.685000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 13.4438 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 66.983 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 68.4163 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 340.88 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 446.635000 0.000000 446.775000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430000 0.000000 933.570000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.520000 0.000000 931.660000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.615000 0.000000 929.755000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.705000 0.000000 927.845000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.795000 0.000000 925.935000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.885000 0.000000 924.025000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.975000 0.000000 922.115000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.070000 0.000000 920.210000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.160000 0.000000 918.300000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.250000 0.000000 916.390000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.340000 0.000000 914.480000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.430000 0.000000 912.570000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.525000 0.000000 910.665000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.615000 0.000000 908.755000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.705000 0.000000 906.845000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.795000 0.000000 904.935000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.885000 0.000000 903.025000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.980000 0.000000 901.120000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.070000 0.000000 899.210000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.160000 0.000000 897.300000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.250000 0.000000 895.390000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.340000 0.000000 893.480000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.435000 0.000000 891.575000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.525000 0.000000 889.665000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.615000 0.000000 887.755000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.705000 0.000000 885.845000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.795000 0.000000 883.935000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.890000 0.000000 882.030000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.980000 0.000000 880.120000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.070000 0.000000 878.210000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.160000 0.000000 876.300000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.250000 0.000000 874.390000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.345000 0.000000 872.485000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.435000 0.000000 870.575000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.525000 0.000000 868.665000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.615000 0.000000 866.755000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.705000 0.000000 864.845000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.800000 0.000000 862.940000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.890000 0.000000 861.030000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.980000 0.000000 859.120000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.070000 0.000000 857.210000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.160000 0.000000 855.300000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.255000 0.000000 853.395000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.345000 0.000000 851.485000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.435000 0.000000 849.575000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.525000 0.000000 847.665000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.615000 0.000000 845.755000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.710000 0.000000 843.850000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.800000 0.000000 841.940000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.890000 0.000000 840.030000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.980000 0.000000 838.120000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.070000 0.000000 836.210000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.165000 0.000000 834.305000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.255000 0.000000 832.395000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.345000 0.000000 830.485000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.435000 0.000000 828.575000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.525000 0.000000 826.665000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.620000 0.000000 824.760000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.710000 0.000000 822.850000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.800000 0.000000 820.940000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890000 0.000000 819.030000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.980000 0.000000 817.120000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1799 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.7385 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 50.6845 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 270.784 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 113.581 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 606.704 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 12.87 LAYER met4  ;
    ANTENNAMAXAREACAR 12.075 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 62.8933 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.0663636 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 815.075000 0.000000 815.215000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7182 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.43 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.231 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 39.032 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 468.024 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2505.03 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 19.056 LAYER met4  ;
    ANTENNAMAXAREACAR 88.5373 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 467.863 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.472525 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 813.165000 0.000000 813.305000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5624 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.651 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.4648 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 13.616 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met3  ;
    ANTENNAMAXAREACAR 13.9774 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 70.9374 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.369293 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 811.255000 0.000000 811.395000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9485 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.5165 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.9034 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 48.004 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 809.345000 0.000000 809.485000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7735 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.6415 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.30707 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.0687 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 807.435000 0.000000 807.575000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.036 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.954 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 13.2707 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 59.8404 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 805.530000 0.000000 805.670000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8101 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.9425 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.63768 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.0222 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 803.620000 0.000000 803.760000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.701 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4501 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 51.2141 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 801.710000 0.000000 801.850000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6498 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.141 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 10.84 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 49.1455 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 799.800000 0.000000 799.940000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.847 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.009 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.4077 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 53.299 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 797.890000 0.000000 798.030000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6043 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.9135 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.57455 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 37.8182 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 795.985000 0.000000 796.125000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0824 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.5185 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 52.4263 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 794.075000 0.000000 794.215000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7149 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4665 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 15.0302 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 71.4008 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 792.165000 0.000000 792.305000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6603 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.1935 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 18.0167 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 80.5556 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 790.255000 0.000000 790.395000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.904 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.14667 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.0586 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 788.345000 0.000000 788.485000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.526 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.30111 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.3394 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 786.440000 0.000000 786.580000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7394 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.589 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.53818 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.6545 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 784.530000 0.000000 784.670000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6988 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.386 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.19737 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.8343 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 782.620000 0.000000 782.760000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6918 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.351 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.4199 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 41.9333 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 780.710000 0.000000 780.850000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7268 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.526 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.1225 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.4465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 778.800000 0.000000 778.940000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1762 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 10.773 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 11.303 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 50.4788 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 776.895000 0.000000 777.035000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6729 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.2565 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.954 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 85.4841 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 774.985000 0.000000 775.125000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6827 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3055 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.67051 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.4727 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 773.075000 0.000000 773.215000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6925 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3545 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 7.66848 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.6465 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 771.165000 0.000000 771.305000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.801 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.897 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 19.6444 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 88.6944 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 769.255000 0.000000 769.395000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7644 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.596 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.47192 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.6202 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 767.350000 0.000000 767.490000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8344 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.946 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 23.4873 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 106.972 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 765.440000 0.000000 765.580000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7618 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.701 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.88889 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 43.4081 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 763.530000 0.000000 763.670000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6092 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.938 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.62101 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 38.9434 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 761.620000 0.000000 761.760000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.561 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 9.06919 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 40.1798 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 759.710000 0.000000 759.850000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6855 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.3195 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 20.4819 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 87.5238 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 757.805000 0.000000 757.945000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7093 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 8.4385 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 17.4683 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 75.2302 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 755.895000 0.000000 756.035000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5392 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.588 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met2  ;
    ANTENNAMAXAREACAR 27.9984 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 135.706 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.407937 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 753.985000 0.000000 754.125000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8505 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.0265 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 8.33394 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 39.3778 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 752.075000 0.000000 752.215000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.165000 0.000000 750.305000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.260000 0.000000 748.400000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.350000 0.000000 746.490000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.440000 0.000000 744.580000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530000 0.000000 742.670000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.620000 0.000000 740.760000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.715000 0.000000 738.855000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.805000 0.000000 736.945000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.895000 0.000000 735.035000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.985000 0.000000 733.125000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.075000 0.000000 731.215000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.170000 0.000000 729.310000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.260000 0.000000 727.400000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.350000 0.000000 725.490000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.440000 0.000000 723.580000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.530000 0.000000 721.670000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.625000 0.000000 719.765000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.715000 0.000000 717.855000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.805000 0.000000 715.945000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.895000 0.000000 714.035000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.985000 0.000000 712.125000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.080000 0.000000 710.220000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.170000 0.000000 708.310000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.260000 0.000000 706.400000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350000 0.000000 704.490000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.440000 0.000000 702.580000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.535000 0.000000 700.675000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.625000 0.000000 698.765000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.715000 0.000000 696.855000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.805000 0.000000 694.945000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9711 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 9.7475 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.318 LAYER met2  ;
    ANTENNAMAXAREACAR 7.86541 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 36.8113 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.161635 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 692.895000 0.000000 693.035000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.990000 0.000000 691.130000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 45.030000 0.800000 45.330000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 112.795000 0.800000 113.095000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 180.560000 0.800000 180.860000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 248.330000 0.800000 248.630000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 316.095000 0.800000 316.395000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 383.865000 0.800000 384.165000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 451.630000 0.800000 451.930000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 519.395000 0.800000 519.695000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 587.165000 0.800000 587.465000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 654.930000 0.800000 655.230000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 722.700000 0.800000 723.000000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 790.465000 0.800000 790.765000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 858.230000 0.800000 858.530000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 916.070000 0.800000 916.370000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.760000 925.670000 71.900000 926.160000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.505000 925.670000 179.645000 926.160000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.250000 925.670000 287.390000 926.160000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.995000 925.670000 395.135000 926.160000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.740000 925.670000 502.880000 926.160000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.485000 925.670000 610.625000 926.160000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.230000 925.670000 718.370000 926.160000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.975000 925.670000 826.115000 926.160000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.720000 925.670000 913.860000 926.160000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 883.910000 933.800000 884.210000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 820.760000 933.800000 821.060000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 757.615000 933.800000 757.915000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 694.465000 933.800000 694.765000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 631.320000 933.800000 631.620000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 568.175000 933.800000 568.475000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 505.025000 933.800000 505.325000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 441.880000 933.800000 442.180000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 378.730000 933.800000 379.030000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6058 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.159 LAYER met4  ;
    ANTENNAMAXAREACAR 60.1553 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 307.34 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.826415 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 315.585000 933.800000 315.885000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 252.440000 933.800000 252.740000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 189.290000 933.800000 189.590000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 126.145000 933.800000 126.445000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 62.995000 933.800000 63.295000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 933.000000 9.610000 933.800000 9.910000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9221 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 17.472 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 30.350000 0.800000 30.650000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 12.6339 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 67.856 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 90.205000 0.800000 90.505000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 77.4639 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 413.616 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 157.975000 0.800000 158.275000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 125.492 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 669.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 225.740000 0.800000 226.040000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 114.976 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 613.68 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 293.505000 0.800000 293.805000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 128.958 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 687.768 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 2.4978 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 13.792 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 361.275000 0.800000 361.575000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2556 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.688 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 37.4652 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 201.696 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 429.040000 0.800000 429.340000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.7586 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 78.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 33.4326 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 179.248 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 496.810000 0.800000 497.110000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 96.0541 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 512.28 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 52.9908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 283.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 564.575000 0.800000 564.875000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.8206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 67.3824 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 360.784 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 632.340000 0.800000 632.640000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 78.1504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 417.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.6736 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 319.2 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 700.110000 0.800000 700.410000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 75.0439 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 400.696 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 47.2458 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 252.448 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 767.875000 0.800000 768.175000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 66.3949 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 354.568 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 106.3 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 567.872 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 835.645000 0.800000 835.945000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 77.3251 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 412.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 148.087 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 790.736 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 903.410000 0.800000 903.710000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7614 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 58.646 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 52.378 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 279.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 121.855 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 650.832 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 35.845000 925.670000 35.985000 926.160000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.4396 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 37.037 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 29.656 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 158.632 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 140.29 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 749.152 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 143.590000 925.670000 143.730000 926.160000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.199 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 50.834 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 34.831 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 186.232 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 144.937 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 773.936 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 251.335000 925.670000 251.475000 926.160000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 3.6645 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.78 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 160.094 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 854.304 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 359.080000 925.670000 359.220000 926.160000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5666 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.672 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 10.3308 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 55.568 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 466.825000 925.670000 466.965000 926.160000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3259 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 11.3505 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 1.435 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.12 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 42.3528 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 226.352 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 574.570000 925.670000 574.710000 926.160000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3834 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 2.4567 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 12.1555 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 682.315000 925.670000 682.455000 926.160000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7291 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 13.3665 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 68.284 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 364.648 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 40.3398 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 215.616 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 790.060000 925.670000 790.200000 926.160000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4313 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.8775 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 83.98 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 448.36 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.7952 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 38.7798 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 207.296 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 897.805000 925.670000 897.945000 926.160000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9541 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.08 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 151.906 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 811.104 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 904.955000 933.800000 905.255000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 68.4094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 365.312 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 34.9848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 187.056 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 841.810000 933.800000 842.110000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 86.8399 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 463.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 25.6038 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 137.024 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 778.665000 933.800000 778.965000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0059 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 21.1638 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 113.344 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 715.515000 933.800000 715.815000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3834 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.2358 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.728 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 652.370000 933.800000 652.670000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0316 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 16.16 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 53.8566 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 288.176 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 313.431 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 1661.96 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 589.220000 933.800000 589.520000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8881 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.728 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.3406 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 12.4518 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 66.88 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 526.075000 933.800000 526.375000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4986 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.984 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.5156 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 153.024 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 177.262 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 939.109 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 462.930000 933.800000 463.230000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 132.549 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 707.392 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.4455 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 28.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 150.944 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 168.038 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 884.239 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.668702 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 399.780000 933.800000 400.080000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5731 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.048 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 336.635000 933.800000 336.935000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 99.5979 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 531.664 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 273.485000 933.800000 273.785000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4216 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.24 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 210.340000 933.800000 210.640000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3121 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 147.195000 933.800000 147.495000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2161 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.144 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 84.045000 933.800000 84.345000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.7672 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 105.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1244 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.696 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met4  ;
    ANTENNAMAXAREACAR 51.6061 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 247.578 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNAMAXCUTCAR 3.9257 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 101.651 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 344.65 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 20.900000 933.800000 21.200000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9791 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.540000 0.000000 0.840000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0641 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 11 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 67.615000 0.800000 67.915000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7491 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.32 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 135.385000 0.800000 135.685000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5886 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 203.150000 0.800000 203.450000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5346 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 270.920000 0.800000 271.220000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5421 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.216 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 338.685000 0.800000 338.985000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6126 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 406.450000 0.800000 406.750000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6516 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 474.220000 0.800000 474.520000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.408 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 541.985000 0.800000 542.285000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4941 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.96 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 609.755000 0.800000 610.055000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6366 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 8.72 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 677.520000 0.800000 677.820000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2781 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 6.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 745.285000 0.800000 745.585000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4341 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 7.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 813.055000 0.800000 813.355000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.787 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.664 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 880.820000 0.800000 881.120000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.511 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.982 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 10.280000 925.670000 10.420000 926.160000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.5395 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.3885 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.982 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 107.675000 925.670000 107.815000 926.160000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.511 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.982 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 215.420000 925.670000 215.560000 926.160000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.564 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 42.511 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 3.982 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 21.704 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 323.165000 925.670000 323.305000 926.160000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4819 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 7.2485 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 2.1735 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 16.3408 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 88.088 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.421 LAYER met3  ;
    ANTENNAMAXAREACAR 11.1958 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 40.6541 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAMAXCUTCAR 0.125343 LAYER via3  ;
    ANTENNADIFFAREA 2.1735 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 175.287 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 928.96 LAYER met4  ;
    ANTENNAGATEAREA 2.421 LAYER met4  ;
    ANTENNAMAXAREACAR 83.5985 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 424.363 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNAMAXCUTCAR 0.65405 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 133.643 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 521.436 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 430.910000 925.670000 431.050000 926.160000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.824 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.3093 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 538.655000 925.670000 538.795000 926.160000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2266 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.824 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.3093 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 646.400000 925.670000 646.540000 926.160000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2021 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.7015 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.3093 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 754.145000 925.670000 754.285000 926.160000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1923 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 5.5545 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 25.3093 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met2 ;
        RECT 861.890000 925.670000 862.030000 926.160000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.1893 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 917.900000 933.800000 918.200000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.1893 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.656 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 862.860000 933.800000 863.160000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.1143 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 799.710000 933.800000 800.010000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.1143 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 736.565000 933.800000 736.865000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.1143 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 137.256 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 673.420000 933.800000 673.720000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.0693 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.536 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.2138 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 8.152 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 0.64 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 610.270000 933.800000 610.570000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8071 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.296 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 18.4097 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 90.4 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 547.125000 933.800000 547.425000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2761 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 19.6907 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 97.232 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 483.975000 933.800000 484.275000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2356 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.248 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 420.830000 933.800000 421.130000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.3365 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.7057 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 341.176 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.3365 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 18.9516 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 102.016 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 9.822 LAYER met4  ;
    ANTENNAMAXAREACAR 35.5207 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 181.959 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.504894 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 357.685000 933.800000 357.985000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4261 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 294.535000 933.800000 294.835000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3166 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 231.390000 933.800000 231.690000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2206 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 168.240000 933.800000 168.540000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3091 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.64 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 105.095000 933.800000 105.395000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2146 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 119.732 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 629.736 LAYER met4  ;
    ANTENNAPARTIALCUTAREA 1.28 LAYER via4  ;
    ANTENNADIFFAREA 2.1735 LAYER met5  ;
    ANTENNAPARTIALMETALAREA 130.992 LAYER met5  ;
    ANTENNAPARTIALMETALSIDEAREA 254.088 LAYER met5  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.6175 LAYER met5  ;
    ANTENNAMAXAREACAR 50.0447 LAYER met5  ;
    ANTENNAMAXSIDEAREACAR 97.0728 LAYER met5  ;
    PORT
      LAYER met3 ;
        RECT 933.000000 41.950000 933.800000 42.250000 ;
    END
  END io_oeb[0]
  PIN irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0421 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 8.390000 0.800000 8.690000 ;
    END
  END irq[2]
  PIN irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0421 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 16.320000 0.800000 16.620000 ;
    END
  END irq[1]
  PIN irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0421 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 18.592 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 257.848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1375.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 24.250000 0.800000 24.550000 ;
    END
  END irq[0]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 929.740000 2.100000 931.740000 924.060000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.060000 2.100000 4.060000 924.060000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 916.385000 516.980000 918.125000 911.760000 ;
      LAYER met4 ;
        RECT 441.065000 516.980000 442.805000 911.760000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 925.740000 6.100000 927.740000 920.060000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.060000 6.100000 8.060000 920.060000 ;
    END

# P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'
    PORT
      LAYER met4 ;
        RECT 444.465000 520.380000 446.205000 908.360000 ;
      LAYER met4 ;
        RECT 912.985000 520.380000 914.725000 908.360000 ;
    END
# end of P/G pin shape extracted from block 'sky130_sram_1kbyte_1rw1r_32x256_8'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 933.800000 926.160000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 933.800000 926.160000 ;
    LAYER met2 ;
      RECT 914.000000 925.530000 933.800000 926.160000 ;
      RECT 898.085000 925.530000 913.580000 926.160000 ;
      RECT 862.170000 925.530000 897.665000 926.160000 ;
      RECT 826.255000 925.530000 861.750000 926.160000 ;
      RECT 790.340000 925.530000 825.835000 926.160000 ;
      RECT 754.425000 925.530000 789.920000 926.160000 ;
      RECT 718.510000 925.530000 754.005000 926.160000 ;
      RECT 682.595000 925.530000 718.090000 926.160000 ;
      RECT 646.680000 925.530000 682.175000 926.160000 ;
      RECT 610.765000 925.530000 646.260000 926.160000 ;
      RECT 574.850000 925.530000 610.345000 926.160000 ;
      RECT 538.935000 925.530000 574.430000 926.160000 ;
      RECT 503.020000 925.530000 538.515000 926.160000 ;
      RECT 467.105000 925.530000 502.600000 926.160000 ;
      RECT 431.190000 925.530000 466.685000 926.160000 ;
      RECT 395.275000 925.530000 430.770000 926.160000 ;
      RECT 359.360000 925.530000 394.855000 926.160000 ;
      RECT 323.445000 925.530000 358.940000 926.160000 ;
      RECT 287.530000 925.530000 323.025000 926.160000 ;
      RECT 251.615000 925.530000 287.110000 926.160000 ;
      RECT 215.700000 925.530000 251.195000 926.160000 ;
      RECT 179.785000 925.530000 215.280000 926.160000 ;
      RECT 143.870000 925.530000 179.365000 926.160000 ;
      RECT 107.955000 925.530000 143.450000 926.160000 ;
      RECT 72.040000 925.530000 107.535000 926.160000 ;
      RECT 36.125000 925.530000 71.620000 926.160000 ;
      RECT 10.560000 925.530000 35.705000 926.160000 ;
      RECT 0.000000 925.530000 10.140000 926.160000 ;
      RECT 0.000000 5.480000 933.800000 925.530000 ;
      RECT 0.630000 5.060000 933.800000 5.480000 ;
      RECT 0.000000 0.630000 933.800000 5.060000 ;
      RECT 933.710000 0.000000 933.800000 0.630000 ;
      RECT 931.800000 0.000000 933.290000 0.630000 ;
      RECT 929.895000 0.000000 931.380000 0.630000 ;
      RECT 927.985000 0.000000 929.475000 0.630000 ;
      RECT 926.075000 0.000000 927.565000 0.630000 ;
      RECT 924.165000 0.000000 925.655000 0.630000 ;
      RECT 922.255000 0.000000 923.745000 0.630000 ;
      RECT 920.350000 0.000000 921.835000 0.630000 ;
      RECT 918.440000 0.000000 919.930000 0.630000 ;
      RECT 916.530000 0.000000 918.020000 0.630000 ;
      RECT 914.620000 0.000000 916.110000 0.630000 ;
      RECT 912.710000 0.000000 914.200000 0.630000 ;
      RECT 910.805000 0.000000 912.290000 0.630000 ;
      RECT 908.895000 0.000000 910.385000 0.630000 ;
      RECT 906.985000 0.000000 908.475000 0.630000 ;
      RECT 905.075000 0.000000 906.565000 0.630000 ;
      RECT 903.165000 0.000000 904.655000 0.630000 ;
      RECT 901.260000 0.000000 902.745000 0.630000 ;
      RECT 899.350000 0.000000 900.840000 0.630000 ;
      RECT 897.440000 0.000000 898.930000 0.630000 ;
      RECT 895.530000 0.000000 897.020000 0.630000 ;
      RECT 893.620000 0.000000 895.110000 0.630000 ;
      RECT 891.715000 0.000000 893.200000 0.630000 ;
      RECT 889.805000 0.000000 891.295000 0.630000 ;
      RECT 887.895000 0.000000 889.385000 0.630000 ;
      RECT 885.985000 0.000000 887.475000 0.630000 ;
      RECT 884.075000 0.000000 885.565000 0.630000 ;
      RECT 882.170000 0.000000 883.655000 0.630000 ;
      RECT 880.260000 0.000000 881.750000 0.630000 ;
      RECT 878.350000 0.000000 879.840000 0.630000 ;
      RECT 876.440000 0.000000 877.930000 0.630000 ;
      RECT 874.530000 0.000000 876.020000 0.630000 ;
      RECT 872.625000 0.000000 874.110000 0.630000 ;
      RECT 870.715000 0.000000 872.205000 0.630000 ;
      RECT 868.805000 0.000000 870.295000 0.630000 ;
      RECT 866.895000 0.000000 868.385000 0.630000 ;
      RECT 864.985000 0.000000 866.475000 0.630000 ;
      RECT 863.080000 0.000000 864.565000 0.630000 ;
      RECT 861.170000 0.000000 862.660000 0.630000 ;
      RECT 859.260000 0.000000 860.750000 0.630000 ;
      RECT 857.350000 0.000000 858.840000 0.630000 ;
      RECT 855.440000 0.000000 856.930000 0.630000 ;
      RECT 853.535000 0.000000 855.020000 0.630000 ;
      RECT 851.625000 0.000000 853.115000 0.630000 ;
      RECT 849.715000 0.000000 851.205000 0.630000 ;
      RECT 847.805000 0.000000 849.295000 0.630000 ;
      RECT 845.895000 0.000000 847.385000 0.630000 ;
      RECT 843.990000 0.000000 845.475000 0.630000 ;
      RECT 842.080000 0.000000 843.570000 0.630000 ;
      RECT 840.170000 0.000000 841.660000 0.630000 ;
      RECT 838.260000 0.000000 839.750000 0.630000 ;
      RECT 836.350000 0.000000 837.840000 0.630000 ;
      RECT 834.445000 0.000000 835.930000 0.630000 ;
      RECT 832.535000 0.000000 834.025000 0.630000 ;
      RECT 830.625000 0.000000 832.115000 0.630000 ;
      RECT 828.715000 0.000000 830.205000 0.630000 ;
      RECT 826.805000 0.000000 828.295000 0.630000 ;
      RECT 824.900000 0.000000 826.385000 0.630000 ;
      RECT 822.990000 0.000000 824.480000 0.630000 ;
      RECT 821.080000 0.000000 822.570000 0.630000 ;
      RECT 819.170000 0.000000 820.660000 0.630000 ;
      RECT 817.260000 0.000000 818.750000 0.630000 ;
      RECT 815.355000 0.000000 816.840000 0.630000 ;
      RECT 813.445000 0.000000 814.935000 0.630000 ;
      RECT 811.535000 0.000000 813.025000 0.630000 ;
      RECT 809.625000 0.000000 811.115000 0.630000 ;
      RECT 807.715000 0.000000 809.205000 0.630000 ;
      RECT 805.810000 0.000000 807.295000 0.630000 ;
      RECT 803.900000 0.000000 805.390000 0.630000 ;
      RECT 801.990000 0.000000 803.480000 0.630000 ;
      RECT 800.080000 0.000000 801.570000 0.630000 ;
      RECT 798.170000 0.000000 799.660000 0.630000 ;
      RECT 796.265000 0.000000 797.750000 0.630000 ;
      RECT 794.355000 0.000000 795.845000 0.630000 ;
      RECT 792.445000 0.000000 793.935000 0.630000 ;
      RECT 790.535000 0.000000 792.025000 0.630000 ;
      RECT 788.625000 0.000000 790.115000 0.630000 ;
      RECT 786.720000 0.000000 788.205000 0.630000 ;
      RECT 784.810000 0.000000 786.300000 0.630000 ;
      RECT 782.900000 0.000000 784.390000 0.630000 ;
      RECT 780.990000 0.000000 782.480000 0.630000 ;
      RECT 779.080000 0.000000 780.570000 0.630000 ;
      RECT 777.175000 0.000000 778.660000 0.630000 ;
      RECT 775.265000 0.000000 776.755000 0.630000 ;
      RECT 773.355000 0.000000 774.845000 0.630000 ;
      RECT 771.445000 0.000000 772.935000 0.630000 ;
      RECT 769.535000 0.000000 771.025000 0.630000 ;
      RECT 767.630000 0.000000 769.115000 0.630000 ;
      RECT 765.720000 0.000000 767.210000 0.630000 ;
      RECT 763.810000 0.000000 765.300000 0.630000 ;
      RECT 761.900000 0.000000 763.390000 0.630000 ;
      RECT 759.990000 0.000000 761.480000 0.630000 ;
      RECT 758.085000 0.000000 759.570000 0.630000 ;
      RECT 756.175000 0.000000 757.665000 0.630000 ;
      RECT 754.265000 0.000000 755.755000 0.630000 ;
      RECT 752.355000 0.000000 753.845000 0.630000 ;
      RECT 750.445000 0.000000 751.935000 0.630000 ;
      RECT 748.540000 0.000000 750.025000 0.630000 ;
      RECT 746.630000 0.000000 748.120000 0.630000 ;
      RECT 744.720000 0.000000 746.210000 0.630000 ;
      RECT 742.810000 0.000000 744.300000 0.630000 ;
      RECT 740.900000 0.000000 742.390000 0.630000 ;
      RECT 738.995000 0.000000 740.480000 0.630000 ;
      RECT 737.085000 0.000000 738.575000 0.630000 ;
      RECT 735.175000 0.000000 736.665000 0.630000 ;
      RECT 733.265000 0.000000 734.755000 0.630000 ;
      RECT 731.355000 0.000000 732.845000 0.630000 ;
      RECT 729.450000 0.000000 730.935000 0.630000 ;
      RECT 727.540000 0.000000 729.030000 0.630000 ;
      RECT 725.630000 0.000000 727.120000 0.630000 ;
      RECT 723.720000 0.000000 725.210000 0.630000 ;
      RECT 721.810000 0.000000 723.300000 0.630000 ;
      RECT 719.905000 0.000000 721.390000 0.630000 ;
      RECT 717.995000 0.000000 719.485000 0.630000 ;
      RECT 716.085000 0.000000 717.575000 0.630000 ;
      RECT 714.175000 0.000000 715.665000 0.630000 ;
      RECT 712.265000 0.000000 713.755000 0.630000 ;
      RECT 710.360000 0.000000 711.845000 0.630000 ;
      RECT 708.450000 0.000000 709.940000 0.630000 ;
      RECT 706.540000 0.000000 708.030000 0.630000 ;
      RECT 704.630000 0.000000 706.120000 0.630000 ;
      RECT 702.720000 0.000000 704.210000 0.630000 ;
      RECT 700.815000 0.000000 702.300000 0.630000 ;
      RECT 698.905000 0.000000 700.395000 0.630000 ;
      RECT 696.995000 0.000000 698.485000 0.630000 ;
      RECT 695.085000 0.000000 696.575000 0.630000 ;
      RECT 693.175000 0.000000 694.665000 0.630000 ;
      RECT 691.270000 0.000000 692.755000 0.630000 ;
      RECT 689.360000 0.000000 690.850000 0.630000 ;
      RECT 687.450000 0.000000 688.940000 0.630000 ;
      RECT 685.540000 0.000000 687.030000 0.630000 ;
      RECT 683.630000 0.000000 685.120000 0.630000 ;
      RECT 681.725000 0.000000 683.210000 0.630000 ;
      RECT 679.815000 0.000000 681.305000 0.630000 ;
      RECT 677.905000 0.000000 679.395000 0.630000 ;
      RECT 675.995000 0.000000 677.485000 0.630000 ;
      RECT 674.085000 0.000000 675.575000 0.630000 ;
      RECT 672.180000 0.000000 673.665000 0.630000 ;
      RECT 670.270000 0.000000 671.760000 0.630000 ;
      RECT 668.360000 0.000000 669.850000 0.630000 ;
      RECT 666.450000 0.000000 667.940000 0.630000 ;
      RECT 664.540000 0.000000 666.030000 0.630000 ;
      RECT 662.635000 0.000000 664.120000 0.630000 ;
      RECT 660.725000 0.000000 662.215000 0.630000 ;
      RECT 658.815000 0.000000 660.305000 0.630000 ;
      RECT 656.905000 0.000000 658.395000 0.630000 ;
      RECT 654.995000 0.000000 656.485000 0.630000 ;
      RECT 653.090000 0.000000 654.575000 0.630000 ;
      RECT 651.180000 0.000000 652.670000 0.630000 ;
      RECT 649.270000 0.000000 650.760000 0.630000 ;
      RECT 647.360000 0.000000 648.850000 0.630000 ;
      RECT 645.450000 0.000000 646.940000 0.630000 ;
      RECT 643.545000 0.000000 645.030000 0.630000 ;
      RECT 641.635000 0.000000 643.125000 0.630000 ;
      RECT 639.725000 0.000000 641.215000 0.630000 ;
      RECT 637.815000 0.000000 639.305000 0.630000 ;
      RECT 635.905000 0.000000 637.395000 0.630000 ;
      RECT 634.000000 0.000000 635.485000 0.630000 ;
      RECT 632.090000 0.000000 633.580000 0.630000 ;
      RECT 630.180000 0.000000 631.670000 0.630000 ;
      RECT 628.270000 0.000000 629.760000 0.630000 ;
      RECT 626.360000 0.000000 627.850000 0.630000 ;
      RECT 624.455000 0.000000 625.940000 0.630000 ;
      RECT 622.545000 0.000000 624.035000 0.630000 ;
      RECT 620.635000 0.000000 622.125000 0.630000 ;
      RECT 618.725000 0.000000 620.215000 0.630000 ;
      RECT 616.815000 0.000000 618.305000 0.630000 ;
      RECT 614.910000 0.000000 616.395000 0.630000 ;
      RECT 613.000000 0.000000 614.490000 0.630000 ;
      RECT 611.090000 0.000000 612.580000 0.630000 ;
      RECT 609.180000 0.000000 610.670000 0.630000 ;
      RECT 607.270000 0.000000 608.760000 0.630000 ;
      RECT 605.365000 0.000000 606.850000 0.630000 ;
      RECT 603.455000 0.000000 604.945000 0.630000 ;
      RECT 601.545000 0.000000 603.035000 0.630000 ;
      RECT 599.635000 0.000000 601.125000 0.630000 ;
      RECT 597.725000 0.000000 599.215000 0.630000 ;
      RECT 595.820000 0.000000 597.305000 0.630000 ;
      RECT 593.910000 0.000000 595.400000 0.630000 ;
      RECT 592.000000 0.000000 593.490000 0.630000 ;
      RECT 590.090000 0.000000 591.580000 0.630000 ;
      RECT 588.180000 0.000000 589.670000 0.630000 ;
      RECT 586.275000 0.000000 587.760000 0.630000 ;
      RECT 584.365000 0.000000 585.855000 0.630000 ;
      RECT 582.455000 0.000000 583.945000 0.630000 ;
      RECT 580.545000 0.000000 582.035000 0.630000 ;
      RECT 578.635000 0.000000 580.125000 0.630000 ;
      RECT 576.730000 0.000000 578.215000 0.630000 ;
      RECT 574.820000 0.000000 576.310000 0.630000 ;
      RECT 572.910000 0.000000 574.400000 0.630000 ;
      RECT 571.000000 0.000000 572.490000 0.630000 ;
      RECT 569.090000 0.000000 570.580000 0.630000 ;
      RECT 567.185000 0.000000 568.670000 0.630000 ;
      RECT 565.275000 0.000000 566.765000 0.630000 ;
      RECT 563.365000 0.000000 564.855000 0.630000 ;
      RECT 561.455000 0.000000 562.945000 0.630000 ;
      RECT 559.545000 0.000000 561.035000 0.630000 ;
      RECT 557.640000 0.000000 559.125000 0.630000 ;
      RECT 555.730000 0.000000 557.220000 0.630000 ;
      RECT 553.820000 0.000000 555.310000 0.630000 ;
      RECT 551.910000 0.000000 553.400000 0.630000 ;
      RECT 550.000000 0.000000 551.490000 0.630000 ;
      RECT 548.095000 0.000000 549.580000 0.630000 ;
      RECT 546.185000 0.000000 547.675000 0.630000 ;
      RECT 544.275000 0.000000 545.765000 0.630000 ;
      RECT 542.365000 0.000000 543.855000 0.630000 ;
      RECT 540.455000 0.000000 541.945000 0.630000 ;
      RECT 538.550000 0.000000 540.035000 0.630000 ;
      RECT 536.640000 0.000000 538.130000 0.630000 ;
      RECT 534.730000 0.000000 536.220000 0.630000 ;
      RECT 532.820000 0.000000 534.310000 0.630000 ;
      RECT 530.910000 0.000000 532.400000 0.630000 ;
      RECT 529.005000 0.000000 530.490000 0.630000 ;
      RECT 527.095000 0.000000 528.585000 0.630000 ;
      RECT 525.185000 0.000000 526.675000 0.630000 ;
      RECT 523.275000 0.000000 524.765000 0.630000 ;
      RECT 521.365000 0.000000 522.855000 0.630000 ;
      RECT 519.460000 0.000000 520.945000 0.630000 ;
      RECT 517.550000 0.000000 519.040000 0.630000 ;
      RECT 515.640000 0.000000 517.130000 0.630000 ;
      RECT 513.730000 0.000000 515.220000 0.630000 ;
      RECT 511.820000 0.000000 513.310000 0.630000 ;
      RECT 509.915000 0.000000 511.400000 0.630000 ;
      RECT 508.005000 0.000000 509.495000 0.630000 ;
      RECT 506.095000 0.000000 507.585000 0.630000 ;
      RECT 504.185000 0.000000 505.675000 0.630000 ;
      RECT 502.275000 0.000000 503.765000 0.630000 ;
      RECT 500.370000 0.000000 501.855000 0.630000 ;
      RECT 498.460000 0.000000 499.950000 0.630000 ;
      RECT 496.550000 0.000000 498.040000 0.630000 ;
      RECT 494.640000 0.000000 496.130000 0.630000 ;
      RECT 492.730000 0.000000 494.220000 0.630000 ;
      RECT 490.825000 0.000000 492.310000 0.630000 ;
      RECT 488.915000 0.000000 490.405000 0.630000 ;
      RECT 487.005000 0.000000 488.495000 0.630000 ;
      RECT 485.095000 0.000000 486.585000 0.630000 ;
      RECT 483.185000 0.000000 484.675000 0.630000 ;
      RECT 481.280000 0.000000 482.765000 0.630000 ;
      RECT 479.370000 0.000000 480.860000 0.630000 ;
      RECT 477.460000 0.000000 478.950000 0.630000 ;
      RECT 475.550000 0.000000 477.040000 0.630000 ;
      RECT 473.640000 0.000000 475.130000 0.630000 ;
      RECT 471.735000 0.000000 473.220000 0.630000 ;
      RECT 469.825000 0.000000 471.315000 0.630000 ;
      RECT 467.915000 0.000000 469.405000 0.630000 ;
      RECT 466.005000 0.000000 467.495000 0.630000 ;
      RECT 464.095000 0.000000 465.585000 0.630000 ;
      RECT 462.190000 0.000000 463.675000 0.630000 ;
      RECT 460.280000 0.000000 461.770000 0.630000 ;
      RECT 458.370000 0.000000 459.860000 0.630000 ;
      RECT 456.460000 0.000000 457.950000 0.630000 ;
      RECT 454.550000 0.000000 456.040000 0.630000 ;
      RECT 452.645000 0.000000 454.130000 0.630000 ;
      RECT 450.735000 0.000000 452.225000 0.630000 ;
      RECT 448.825000 0.000000 450.315000 0.630000 ;
      RECT 446.915000 0.000000 448.405000 0.630000 ;
      RECT 445.005000 0.000000 446.495000 0.630000 ;
      RECT 443.100000 0.000000 444.585000 0.630000 ;
      RECT 441.190000 0.000000 442.680000 0.630000 ;
      RECT 439.280000 0.000000 440.770000 0.630000 ;
      RECT 437.370000 0.000000 438.860000 0.630000 ;
      RECT 435.460000 0.000000 436.950000 0.630000 ;
      RECT 433.555000 0.000000 435.040000 0.630000 ;
      RECT 431.645000 0.000000 433.135000 0.630000 ;
      RECT 429.735000 0.000000 431.225000 0.630000 ;
      RECT 427.825000 0.000000 429.315000 0.630000 ;
      RECT 425.915000 0.000000 427.405000 0.630000 ;
      RECT 424.010000 0.000000 425.495000 0.630000 ;
      RECT 422.100000 0.000000 423.590000 0.630000 ;
      RECT 420.190000 0.000000 421.680000 0.630000 ;
      RECT 418.280000 0.000000 419.770000 0.630000 ;
      RECT 416.370000 0.000000 417.860000 0.630000 ;
      RECT 414.465000 0.000000 415.950000 0.630000 ;
      RECT 412.555000 0.000000 414.045000 0.630000 ;
      RECT 410.645000 0.000000 412.135000 0.630000 ;
      RECT 408.735000 0.000000 410.225000 0.630000 ;
      RECT 406.825000 0.000000 408.315000 0.630000 ;
      RECT 404.920000 0.000000 406.405000 0.630000 ;
      RECT 403.010000 0.000000 404.500000 0.630000 ;
      RECT 401.100000 0.000000 402.590000 0.630000 ;
      RECT 399.190000 0.000000 400.680000 0.630000 ;
      RECT 397.280000 0.000000 398.770000 0.630000 ;
      RECT 395.375000 0.000000 396.860000 0.630000 ;
      RECT 393.465000 0.000000 394.955000 0.630000 ;
      RECT 391.555000 0.000000 393.045000 0.630000 ;
      RECT 389.645000 0.000000 391.135000 0.630000 ;
      RECT 387.735000 0.000000 389.225000 0.630000 ;
      RECT 385.830000 0.000000 387.315000 0.630000 ;
      RECT 383.920000 0.000000 385.410000 0.630000 ;
      RECT 382.010000 0.000000 383.500000 0.630000 ;
      RECT 380.100000 0.000000 381.590000 0.630000 ;
      RECT 378.190000 0.000000 379.680000 0.630000 ;
      RECT 376.285000 0.000000 377.770000 0.630000 ;
      RECT 374.375000 0.000000 375.865000 0.630000 ;
      RECT 372.465000 0.000000 373.955000 0.630000 ;
      RECT 370.555000 0.000000 372.045000 0.630000 ;
      RECT 368.645000 0.000000 370.135000 0.630000 ;
      RECT 366.740000 0.000000 368.225000 0.630000 ;
      RECT 364.830000 0.000000 366.320000 0.630000 ;
      RECT 362.920000 0.000000 364.410000 0.630000 ;
      RECT 361.010000 0.000000 362.500000 0.630000 ;
      RECT 359.100000 0.000000 360.590000 0.630000 ;
      RECT 357.195000 0.000000 358.680000 0.630000 ;
      RECT 355.285000 0.000000 356.775000 0.630000 ;
      RECT 353.375000 0.000000 354.865000 0.630000 ;
      RECT 351.465000 0.000000 352.955000 0.630000 ;
      RECT 349.555000 0.000000 351.045000 0.630000 ;
      RECT 347.650000 0.000000 349.135000 0.630000 ;
      RECT 345.740000 0.000000 347.230000 0.630000 ;
      RECT 343.830000 0.000000 345.320000 0.630000 ;
      RECT 341.920000 0.000000 343.410000 0.630000 ;
      RECT 340.010000 0.000000 341.500000 0.630000 ;
      RECT 338.105000 0.000000 339.590000 0.630000 ;
      RECT 336.195000 0.000000 337.685000 0.630000 ;
      RECT 334.285000 0.000000 335.775000 0.630000 ;
      RECT 332.375000 0.000000 333.865000 0.630000 ;
      RECT 330.465000 0.000000 331.955000 0.630000 ;
      RECT 328.560000 0.000000 330.045000 0.630000 ;
      RECT 326.650000 0.000000 328.140000 0.630000 ;
      RECT 324.740000 0.000000 326.230000 0.630000 ;
      RECT 322.830000 0.000000 324.320000 0.630000 ;
      RECT 320.920000 0.000000 322.410000 0.630000 ;
      RECT 319.015000 0.000000 320.500000 0.630000 ;
      RECT 317.105000 0.000000 318.595000 0.630000 ;
      RECT 315.195000 0.000000 316.685000 0.630000 ;
      RECT 313.285000 0.000000 314.775000 0.630000 ;
      RECT 311.375000 0.000000 312.865000 0.630000 ;
      RECT 309.470000 0.000000 310.955000 0.630000 ;
      RECT 307.560000 0.000000 309.050000 0.630000 ;
      RECT 305.650000 0.000000 307.140000 0.630000 ;
      RECT 303.740000 0.000000 305.230000 0.630000 ;
      RECT 301.830000 0.000000 303.320000 0.630000 ;
      RECT 299.925000 0.000000 301.410000 0.630000 ;
      RECT 298.015000 0.000000 299.505000 0.630000 ;
      RECT 296.105000 0.000000 297.595000 0.630000 ;
      RECT 294.195000 0.000000 295.685000 0.630000 ;
      RECT 292.285000 0.000000 293.775000 0.630000 ;
      RECT 290.380000 0.000000 291.865000 0.630000 ;
      RECT 288.470000 0.000000 289.960000 0.630000 ;
      RECT 286.560000 0.000000 288.050000 0.630000 ;
      RECT 284.650000 0.000000 286.140000 0.630000 ;
      RECT 282.740000 0.000000 284.230000 0.630000 ;
      RECT 280.835000 0.000000 282.320000 0.630000 ;
      RECT 278.925000 0.000000 280.415000 0.630000 ;
      RECT 277.015000 0.000000 278.505000 0.630000 ;
      RECT 275.105000 0.000000 276.595000 0.630000 ;
      RECT 273.195000 0.000000 274.685000 0.630000 ;
      RECT 271.290000 0.000000 272.775000 0.630000 ;
      RECT 269.380000 0.000000 270.870000 0.630000 ;
      RECT 267.470000 0.000000 268.960000 0.630000 ;
      RECT 265.560000 0.000000 267.050000 0.630000 ;
      RECT 263.650000 0.000000 265.140000 0.630000 ;
      RECT 261.745000 0.000000 263.230000 0.630000 ;
      RECT 259.835000 0.000000 261.325000 0.630000 ;
      RECT 257.925000 0.000000 259.415000 0.630000 ;
      RECT 256.015000 0.000000 257.505000 0.630000 ;
      RECT 254.105000 0.000000 255.595000 0.630000 ;
      RECT 252.200000 0.000000 253.685000 0.630000 ;
      RECT 250.290000 0.000000 251.780000 0.630000 ;
      RECT 248.380000 0.000000 249.870000 0.630000 ;
      RECT 246.470000 0.000000 247.960000 0.630000 ;
      RECT 244.560000 0.000000 246.050000 0.630000 ;
      RECT 242.655000 0.000000 244.140000 0.630000 ;
      RECT 240.745000 0.000000 242.235000 0.630000 ;
      RECT 238.835000 0.000000 240.325000 0.630000 ;
      RECT 236.925000 0.000000 238.415000 0.630000 ;
      RECT 235.015000 0.000000 236.505000 0.630000 ;
      RECT 233.110000 0.000000 234.595000 0.630000 ;
      RECT 231.200000 0.000000 232.690000 0.630000 ;
      RECT 229.290000 0.000000 230.780000 0.630000 ;
      RECT 227.380000 0.000000 228.870000 0.630000 ;
      RECT 225.470000 0.000000 226.960000 0.630000 ;
      RECT 223.565000 0.000000 225.050000 0.630000 ;
      RECT 221.655000 0.000000 223.145000 0.630000 ;
      RECT 219.745000 0.000000 221.235000 0.630000 ;
      RECT 217.835000 0.000000 219.325000 0.630000 ;
      RECT 215.925000 0.000000 217.415000 0.630000 ;
      RECT 214.020000 0.000000 215.505000 0.630000 ;
      RECT 212.110000 0.000000 213.600000 0.630000 ;
      RECT 210.200000 0.000000 211.690000 0.630000 ;
      RECT 208.290000 0.000000 209.780000 0.630000 ;
      RECT 206.380000 0.000000 207.870000 0.630000 ;
      RECT 204.475000 0.000000 205.960000 0.630000 ;
      RECT 202.565000 0.000000 204.055000 0.630000 ;
      RECT 200.655000 0.000000 202.145000 0.630000 ;
      RECT 198.745000 0.000000 200.235000 0.630000 ;
      RECT 196.835000 0.000000 198.325000 0.630000 ;
      RECT 194.930000 0.000000 196.415000 0.630000 ;
      RECT 193.020000 0.000000 194.510000 0.630000 ;
      RECT 191.110000 0.000000 192.600000 0.630000 ;
      RECT 189.200000 0.000000 190.690000 0.630000 ;
      RECT 187.290000 0.000000 188.780000 0.630000 ;
      RECT 185.385000 0.000000 186.870000 0.630000 ;
      RECT 183.475000 0.000000 184.965000 0.630000 ;
      RECT 181.565000 0.000000 183.055000 0.630000 ;
      RECT 179.655000 0.000000 181.145000 0.630000 ;
      RECT 177.745000 0.000000 179.235000 0.630000 ;
      RECT 175.840000 0.000000 177.325000 0.630000 ;
      RECT 173.930000 0.000000 175.420000 0.630000 ;
      RECT 172.020000 0.000000 173.510000 0.630000 ;
      RECT 170.110000 0.000000 171.600000 0.630000 ;
      RECT 168.200000 0.000000 169.690000 0.630000 ;
      RECT 166.295000 0.000000 167.780000 0.630000 ;
      RECT 164.385000 0.000000 165.875000 0.630000 ;
      RECT 162.475000 0.000000 163.965000 0.630000 ;
      RECT 160.565000 0.000000 162.055000 0.630000 ;
      RECT 158.655000 0.000000 160.145000 0.630000 ;
      RECT 156.750000 0.000000 158.235000 0.630000 ;
      RECT 154.840000 0.000000 156.330000 0.630000 ;
      RECT 152.930000 0.000000 154.420000 0.630000 ;
      RECT 151.020000 0.000000 152.510000 0.630000 ;
      RECT 149.110000 0.000000 150.600000 0.630000 ;
      RECT 147.205000 0.000000 148.690000 0.630000 ;
      RECT 145.295000 0.000000 146.785000 0.630000 ;
      RECT 143.385000 0.000000 144.875000 0.630000 ;
      RECT 141.475000 0.000000 142.965000 0.630000 ;
      RECT 139.565000 0.000000 141.055000 0.630000 ;
      RECT 137.660000 0.000000 139.145000 0.630000 ;
      RECT 135.750000 0.000000 137.240000 0.630000 ;
      RECT 133.840000 0.000000 135.330000 0.630000 ;
      RECT 131.930000 0.000000 133.420000 0.630000 ;
      RECT 130.020000 0.000000 131.510000 0.630000 ;
      RECT 128.115000 0.000000 129.600000 0.630000 ;
      RECT 126.205000 0.000000 127.695000 0.630000 ;
      RECT 124.295000 0.000000 125.785000 0.630000 ;
      RECT 122.385000 0.000000 123.875000 0.630000 ;
      RECT 120.475000 0.000000 121.965000 0.630000 ;
      RECT 118.570000 0.000000 120.055000 0.630000 ;
      RECT 116.660000 0.000000 118.150000 0.630000 ;
      RECT 114.750000 0.000000 116.240000 0.630000 ;
      RECT 112.840000 0.000000 114.330000 0.630000 ;
      RECT 110.930000 0.000000 112.420000 0.630000 ;
      RECT 109.025000 0.000000 110.510000 0.630000 ;
      RECT 107.115000 0.000000 108.605000 0.630000 ;
      RECT 105.205000 0.000000 106.695000 0.630000 ;
      RECT 103.295000 0.000000 104.785000 0.630000 ;
      RECT 101.385000 0.000000 102.875000 0.630000 ;
      RECT 99.480000 0.000000 100.965000 0.630000 ;
      RECT 97.570000 0.000000 99.060000 0.630000 ;
      RECT 95.660000 0.000000 97.150000 0.630000 ;
      RECT 93.750000 0.000000 95.240000 0.630000 ;
      RECT 91.840000 0.000000 93.330000 0.630000 ;
      RECT 89.935000 0.000000 91.420000 0.630000 ;
      RECT 88.025000 0.000000 89.515000 0.630000 ;
      RECT 86.115000 0.000000 87.605000 0.630000 ;
      RECT 84.205000 0.000000 85.695000 0.630000 ;
      RECT 82.295000 0.000000 83.785000 0.630000 ;
      RECT 80.390000 0.000000 81.875000 0.630000 ;
      RECT 78.480000 0.000000 79.970000 0.630000 ;
      RECT 76.570000 0.000000 78.060000 0.630000 ;
      RECT 74.660000 0.000000 76.150000 0.630000 ;
      RECT 72.750000 0.000000 74.240000 0.630000 ;
      RECT 70.845000 0.000000 72.330000 0.630000 ;
      RECT 68.935000 0.000000 70.425000 0.630000 ;
      RECT 67.025000 0.000000 68.515000 0.630000 ;
      RECT 65.115000 0.000000 66.605000 0.630000 ;
      RECT 63.205000 0.000000 64.695000 0.630000 ;
      RECT 61.300000 0.000000 62.785000 0.630000 ;
      RECT 59.390000 0.000000 60.880000 0.630000 ;
      RECT 57.480000 0.000000 58.970000 0.630000 ;
      RECT 55.570000 0.000000 57.060000 0.630000 ;
      RECT 53.660000 0.000000 55.150000 0.630000 ;
      RECT 51.755000 0.000000 53.240000 0.630000 ;
      RECT 49.845000 0.000000 51.335000 0.630000 ;
      RECT 47.935000 0.000000 49.425000 0.630000 ;
      RECT 46.025000 0.000000 47.515000 0.630000 ;
      RECT 44.115000 0.000000 45.605000 0.630000 ;
      RECT 42.210000 0.000000 43.695000 0.630000 ;
      RECT 40.300000 0.000000 41.790000 0.630000 ;
      RECT 38.390000 0.000000 39.880000 0.630000 ;
      RECT 36.480000 0.000000 37.970000 0.630000 ;
      RECT 34.570000 0.000000 36.060000 0.630000 ;
      RECT 32.665000 0.000000 34.150000 0.630000 ;
      RECT 30.755000 0.000000 32.245000 0.630000 ;
      RECT 28.845000 0.000000 30.335000 0.630000 ;
      RECT 26.935000 0.000000 28.425000 0.630000 ;
      RECT 25.025000 0.000000 26.515000 0.630000 ;
      RECT 23.120000 0.000000 24.605000 0.630000 ;
      RECT 21.210000 0.000000 22.700000 0.630000 ;
      RECT 19.300000 0.000000 20.790000 0.630000 ;
      RECT 17.390000 0.000000 18.880000 0.630000 ;
      RECT 15.480000 0.000000 16.970000 0.630000 ;
      RECT 13.575000 0.000000 15.060000 0.630000 ;
      RECT 11.665000 0.000000 13.155000 0.630000 ;
      RECT 9.755000 0.000000 11.245000 0.630000 ;
      RECT 7.845000 0.000000 9.335000 0.630000 ;
      RECT 5.935000 0.000000 7.425000 0.630000 ;
      RECT 4.030000 0.000000 5.515000 0.630000 ;
      RECT 2.120000 0.000000 3.610000 0.630000 ;
      RECT 0.000000 0.000000 1.700000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 918.500000 933.800000 926.160000 ;
      RECT 0.000000 917.600000 932.700000 918.500000 ;
      RECT 0.000000 916.670000 933.800000 917.600000 ;
      RECT 1.100000 915.770000 933.800000 916.670000 ;
      RECT 0.000000 905.555000 933.800000 915.770000 ;
      RECT 0.000000 904.655000 932.700000 905.555000 ;
      RECT 0.000000 904.010000 933.800000 904.655000 ;
      RECT 1.100000 903.110000 933.800000 904.010000 ;
      RECT 0.000000 884.510000 933.800000 903.110000 ;
      RECT 0.000000 883.610000 932.700000 884.510000 ;
      RECT 0.000000 881.420000 933.800000 883.610000 ;
      RECT 1.100000 880.520000 933.800000 881.420000 ;
      RECT 0.000000 863.460000 933.800000 880.520000 ;
      RECT 0.000000 862.560000 932.700000 863.460000 ;
      RECT 0.000000 858.830000 933.800000 862.560000 ;
      RECT 1.100000 857.930000 933.800000 858.830000 ;
      RECT 0.000000 842.410000 933.800000 857.930000 ;
      RECT 0.000000 841.510000 932.700000 842.410000 ;
      RECT 0.000000 836.245000 933.800000 841.510000 ;
      RECT 1.100000 835.345000 933.800000 836.245000 ;
      RECT 0.000000 821.360000 933.800000 835.345000 ;
      RECT 0.000000 820.460000 932.700000 821.360000 ;
      RECT 0.000000 813.655000 933.800000 820.460000 ;
      RECT 1.100000 812.755000 933.800000 813.655000 ;
      RECT 0.000000 800.310000 933.800000 812.755000 ;
      RECT 0.000000 799.410000 932.700000 800.310000 ;
      RECT 0.000000 791.065000 933.800000 799.410000 ;
      RECT 1.100000 790.165000 933.800000 791.065000 ;
      RECT 0.000000 779.265000 933.800000 790.165000 ;
      RECT 0.000000 778.365000 932.700000 779.265000 ;
      RECT 0.000000 768.475000 933.800000 778.365000 ;
      RECT 1.100000 767.575000 933.800000 768.475000 ;
      RECT 0.000000 758.215000 933.800000 767.575000 ;
      RECT 0.000000 757.315000 932.700000 758.215000 ;
      RECT 0.000000 745.885000 933.800000 757.315000 ;
      RECT 1.100000 744.985000 933.800000 745.885000 ;
      RECT 0.000000 737.165000 933.800000 744.985000 ;
      RECT 0.000000 736.265000 932.700000 737.165000 ;
      RECT 0.000000 723.300000 933.800000 736.265000 ;
      RECT 1.100000 722.400000 933.800000 723.300000 ;
      RECT 0.000000 716.115000 933.800000 722.400000 ;
      RECT 0.000000 715.215000 932.700000 716.115000 ;
      RECT 0.000000 700.710000 933.800000 715.215000 ;
      RECT 1.100000 699.810000 933.800000 700.710000 ;
      RECT 0.000000 695.065000 933.800000 699.810000 ;
      RECT 0.000000 694.165000 932.700000 695.065000 ;
      RECT 0.000000 678.120000 933.800000 694.165000 ;
      RECT 1.100000 677.220000 933.800000 678.120000 ;
      RECT 0.000000 674.020000 933.800000 677.220000 ;
      RECT 0.000000 673.120000 932.700000 674.020000 ;
      RECT 0.000000 655.530000 933.800000 673.120000 ;
      RECT 1.100000 654.630000 933.800000 655.530000 ;
      RECT 0.000000 652.970000 933.800000 654.630000 ;
      RECT 0.000000 652.070000 932.700000 652.970000 ;
      RECT 0.000000 632.940000 933.800000 652.070000 ;
      RECT 1.100000 632.040000 933.800000 632.940000 ;
      RECT 0.000000 631.920000 933.800000 632.040000 ;
      RECT 0.000000 631.020000 932.700000 631.920000 ;
      RECT 0.000000 610.870000 933.800000 631.020000 ;
      RECT 0.000000 610.355000 932.700000 610.870000 ;
      RECT 1.100000 609.970000 932.700000 610.355000 ;
      RECT 1.100000 609.455000 933.800000 609.970000 ;
      RECT 0.000000 589.820000 933.800000 609.455000 ;
      RECT 0.000000 588.920000 932.700000 589.820000 ;
      RECT 0.000000 587.765000 933.800000 588.920000 ;
      RECT 1.100000 586.865000 933.800000 587.765000 ;
      RECT 0.000000 568.775000 933.800000 586.865000 ;
      RECT 0.000000 567.875000 932.700000 568.775000 ;
      RECT 0.000000 565.175000 933.800000 567.875000 ;
      RECT 1.100000 564.275000 933.800000 565.175000 ;
      RECT 0.000000 547.725000 933.800000 564.275000 ;
      RECT 0.000000 546.825000 932.700000 547.725000 ;
      RECT 0.000000 542.585000 933.800000 546.825000 ;
      RECT 1.100000 541.685000 933.800000 542.585000 ;
      RECT 0.000000 526.675000 933.800000 541.685000 ;
      RECT 0.000000 525.775000 932.700000 526.675000 ;
      RECT 0.000000 519.995000 933.800000 525.775000 ;
      RECT 1.100000 519.095000 933.800000 519.995000 ;
      RECT 0.000000 505.625000 933.800000 519.095000 ;
      RECT 0.000000 504.725000 932.700000 505.625000 ;
      RECT 0.000000 497.410000 933.800000 504.725000 ;
      RECT 1.100000 496.510000 933.800000 497.410000 ;
      RECT 0.000000 484.575000 933.800000 496.510000 ;
      RECT 0.000000 483.675000 932.700000 484.575000 ;
      RECT 0.000000 474.820000 933.800000 483.675000 ;
      RECT 1.100000 473.920000 933.800000 474.820000 ;
      RECT 0.000000 463.530000 933.800000 473.920000 ;
      RECT 0.000000 462.630000 932.700000 463.530000 ;
      RECT 0.000000 452.230000 933.800000 462.630000 ;
      RECT 1.100000 451.330000 933.800000 452.230000 ;
      RECT 0.000000 442.480000 933.800000 451.330000 ;
      RECT 0.000000 441.580000 932.700000 442.480000 ;
      RECT 0.000000 429.640000 933.800000 441.580000 ;
      RECT 1.100000 428.740000 933.800000 429.640000 ;
      RECT 0.000000 421.430000 933.800000 428.740000 ;
      RECT 0.000000 420.530000 932.700000 421.430000 ;
      RECT 0.000000 407.050000 933.800000 420.530000 ;
      RECT 1.100000 406.150000 933.800000 407.050000 ;
      RECT 0.000000 400.380000 933.800000 406.150000 ;
      RECT 0.000000 399.480000 932.700000 400.380000 ;
      RECT 0.000000 384.465000 933.800000 399.480000 ;
      RECT 1.100000 383.565000 933.800000 384.465000 ;
      RECT 0.000000 379.330000 933.800000 383.565000 ;
      RECT 0.000000 378.430000 932.700000 379.330000 ;
      RECT 0.000000 361.875000 933.800000 378.430000 ;
      RECT 1.100000 360.975000 933.800000 361.875000 ;
      RECT 0.000000 358.285000 933.800000 360.975000 ;
      RECT 0.000000 357.385000 932.700000 358.285000 ;
      RECT 0.000000 339.285000 933.800000 357.385000 ;
      RECT 1.100000 338.385000 933.800000 339.285000 ;
      RECT 0.000000 337.235000 933.800000 338.385000 ;
      RECT 0.000000 336.335000 932.700000 337.235000 ;
      RECT 0.000000 316.695000 933.800000 336.335000 ;
      RECT 1.100000 316.185000 933.800000 316.695000 ;
      RECT 1.100000 315.795000 932.700000 316.185000 ;
      RECT 0.000000 315.285000 932.700000 315.795000 ;
      RECT 0.000000 295.135000 933.800000 315.285000 ;
      RECT 0.000000 294.235000 932.700000 295.135000 ;
      RECT 0.000000 294.105000 933.800000 294.235000 ;
      RECT 1.100000 293.205000 933.800000 294.105000 ;
      RECT 0.000000 274.085000 933.800000 293.205000 ;
      RECT 0.000000 273.185000 932.700000 274.085000 ;
      RECT 0.000000 271.520000 933.800000 273.185000 ;
      RECT 1.100000 270.620000 933.800000 271.520000 ;
      RECT 0.000000 253.040000 933.800000 270.620000 ;
      RECT 0.000000 252.140000 932.700000 253.040000 ;
      RECT 0.000000 248.930000 933.800000 252.140000 ;
      RECT 1.100000 248.030000 933.800000 248.930000 ;
      RECT 0.000000 231.990000 933.800000 248.030000 ;
      RECT 0.000000 231.090000 932.700000 231.990000 ;
      RECT 0.000000 226.340000 933.800000 231.090000 ;
      RECT 1.100000 225.440000 933.800000 226.340000 ;
      RECT 0.000000 210.940000 933.800000 225.440000 ;
      RECT 0.000000 210.040000 932.700000 210.940000 ;
      RECT 0.000000 203.750000 933.800000 210.040000 ;
      RECT 1.100000 202.850000 933.800000 203.750000 ;
      RECT 0.000000 189.890000 933.800000 202.850000 ;
      RECT 0.000000 188.990000 932.700000 189.890000 ;
      RECT 0.000000 181.160000 933.800000 188.990000 ;
      RECT 1.100000 180.260000 933.800000 181.160000 ;
      RECT 0.000000 168.840000 933.800000 180.260000 ;
      RECT 0.000000 167.940000 932.700000 168.840000 ;
      RECT 0.000000 158.575000 933.800000 167.940000 ;
      RECT 1.100000 157.675000 933.800000 158.575000 ;
      RECT 0.000000 147.795000 933.800000 157.675000 ;
      RECT 0.000000 146.895000 932.700000 147.795000 ;
      RECT 0.000000 135.985000 933.800000 146.895000 ;
      RECT 1.100000 135.085000 933.800000 135.985000 ;
      RECT 0.000000 126.745000 933.800000 135.085000 ;
      RECT 0.000000 125.845000 932.700000 126.745000 ;
      RECT 0.000000 113.395000 933.800000 125.845000 ;
      RECT 1.100000 112.495000 933.800000 113.395000 ;
      RECT 0.000000 105.695000 933.800000 112.495000 ;
      RECT 0.000000 104.795000 932.700000 105.695000 ;
      RECT 0.000000 90.805000 933.800000 104.795000 ;
      RECT 1.100000 89.905000 933.800000 90.805000 ;
      RECT 0.000000 84.645000 933.800000 89.905000 ;
      RECT 0.000000 83.745000 932.700000 84.645000 ;
      RECT 0.000000 68.215000 933.800000 83.745000 ;
      RECT 1.100000 67.315000 933.800000 68.215000 ;
      RECT 0.000000 63.595000 933.800000 67.315000 ;
      RECT 0.000000 62.695000 932.700000 63.595000 ;
      RECT 0.000000 45.630000 933.800000 62.695000 ;
      RECT 1.100000 44.730000 933.800000 45.630000 ;
      RECT 0.000000 42.550000 933.800000 44.730000 ;
      RECT 0.000000 41.650000 932.700000 42.550000 ;
      RECT 0.000000 30.950000 933.800000 41.650000 ;
      RECT 1.100000 30.050000 933.800000 30.950000 ;
      RECT 0.000000 24.850000 933.800000 30.050000 ;
      RECT 1.100000 23.950000 933.800000 24.850000 ;
      RECT 0.000000 21.500000 933.800000 23.950000 ;
      RECT 0.000000 20.600000 932.700000 21.500000 ;
      RECT 0.000000 16.920000 933.800000 20.600000 ;
      RECT 1.100000 16.020000 933.800000 16.920000 ;
      RECT 0.000000 10.210000 933.800000 16.020000 ;
      RECT 0.000000 9.310000 932.700000 10.210000 ;
      RECT 0.000000 8.990000 933.800000 9.310000 ;
      RECT 1.100000 8.090000 933.800000 8.990000 ;
      RECT 0.000000 1.100000 933.800000 8.090000 ;
      RECT 1.140000 0.000000 933.800000 1.100000 ;
      RECT 0.000000 0.000000 0.240000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 924.360000 933.800000 926.160000 ;
      RECT 4.360000 920.360000 929.440000 924.360000 ;
      RECT 928.040000 5.800000 929.440000 920.360000 ;
      RECT 8.360000 5.800000 925.440000 920.360000 ;
      RECT 4.360000 5.800000 5.760000 920.360000 ;
      RECT 932.040000 1.800000 933.800000 924.360000 ;
      RECT 4.360000 1.800000 929.440000 5.800000 ;
      RECT 0.000000 1.800000 1.760000 924.360000 ;
      RECT 0.000000 0.000000 933.800000 1.800000 ;
  END
END user_proj_example

END LIBRARY
